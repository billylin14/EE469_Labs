//module ARM64BitRegister (clk, ReadRegister1, ReadRegister2, 
//	WriteRegister, WriteData, ReadData1, ReadData2, RegWrite);
//	
//	input logic [4:0] ReadRegister1, ReadRegister2, WriteRegister;
//
//	
//endmodule
	