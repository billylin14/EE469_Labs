module alu (A, B, cntrl, result, negative, zero, overflow, carry_out);

	input logic		[63:0]	A, B;
	input logic		[2:0]		cntrl;
	output logic	[63:0]	result;
	output logic				negative, zero, overflow, carry_out ;
endmodule
